module framer();

endmodule